-------------------------------------------------------------------------------
--
-- Title       : ELEVATOR
-- Design      : ELEVATOR
-- Author      : 
-- Company     : 
--
-------------------------------------------------------------------------------
--
-- File        : ELEVATOR.vhd
-- Generated   : Wed Jul 22 12:01:56 2020
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {ELEVATOR} architecture {ELEVATOR}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

entity ELEVATOR is 
	
	port (
	clk 				:in std_logic; -- clock for the circuit
	ONE_SECOND_CLOCK	:in std_logic; -- clock for counting
	Reset 				:in std_logic;
	start 				:in std_logic;
	
	-- bringing middle signals to the ports to watch them in simulation
	pres_floor			:out std_logic_vector (3 downto 0);	
	targ_floor			:out std_logic_vector (3 downto 0);
	trans_time			:out std_logic_vector (3 downto 0);
	wait_time			:out std_logic_vector (3 downto 0);
	address				:out std_logic_vector (5 downto 0);
	rand_floor			:out std_logic_vector (3 downto 0);
	inter				:out std_logic;
	counter_down		:out integer;
	time_initial		:out integer;
	state				:out std_ulogic_vector(3 downto 0);
	Memory_Out          :out std_logic_vector (7 downto 0);
	
	-- output signals
	Floor 				:out std_logic_vector (3 downto 0);	 
	Timer 				:out std_logic_vector (3 downto 0);
	LiftDir 			:out std_logic_vector (1 downto 0);
	LiftDoor  			:out std_logic	
	);
end ELEVATOR;

--}} End of automatically maintained section

architecture RTL of ELEVATOR is	
-- additional states are present to prevent the compiler from ignoring others (8 states) 
subtype states is std_ulogic_vector(3 downto 0);
constant S0: states 	:= "0000";
constant S1: states 	:= "0001";
constant S2: states 	:= "0010";
constant S3: states 	:= "0011";
constant S4: states 	:= "0100";
constant S5: states 	:= "0101"; 
constant S6: states 	:= "0110";
constant S7: states 	:= "0111";
constant S8: states 	:= "1000";
constant S9: states 	:= "1001"; 
constant S10: states 	:= "1010";
constant S11: states 	:= "1011";
constant S12: states 	:= "1100";
constant S13: states 	:= "1101";
constant S14: states 	:= "1110";
constant finish: states := "1111";

signal fsm_state: std_ulogic_vector(3 downto 0); --for saving the state of the fsm
signal pr_state, nx_state: states;	


-- SOME HELPFUL MIDDLE SIGNALS
signal present_floor 	: std_logic_vector (3 downto 0); -- for saving the current floor
signal target_floor		: std_logic_vector (3 downto 0); -- for saving the target floor	
signal transition_time 	: std_logic_vector (3 downto 0); -- for saving the transition time between two floors
signal waiting_time 	: std_logic_vector (3 downto 0); -- for saving the waiting time of a floor	
signal memory_data 		: std_logic_vector (7 downto 0); -- 8-bit MEMORY data
signal Addr 			: std_logic_vector (5 downto 0); -- 6-bit address  
signal random_floor 	: std_logic_vector (3 downto 0); -- a random floor generated by our LFSR circuit 
signal interrupt 		: std_logic;  -- from random circuit to create interrupt 	 
signal count   			: integer;	  -- for counting the time in the NEXT-STATE-LOGIC process
signal time_init 		: integer range 0 to 20;    -- for initializing the time in seconds, for the COUNTING process


begin 	
	
	
-- S0 : THE STATE BEFORE START HAPPENS FOR INITIALIZATION (WE GO TO THIS STATE WHENEVER RESET IS ON)
-- S1:  FETCHING DATA FROM THE MEMORY
-- S2:  DETERMINES THAT BASED ON THE MEMORY DATA, WE SHOULD GO TO FINISH OR PROCEED TO S3
-- S3:  STATE FOR INITIALIZING time_init WITH TRANSITION TIME
-- S4:  STATE FOR PASSING THE TRANSITION TIME
-- S5:  STATE FOR INITIALIZING time_init WITH WAITING TIME
-- S6:  STATE FOR PASSING WAITING TIME
-- S7:  FROM THIS STATE WE EITHER GO TO S8 FOR A RESPONSE TO INTERRUPT OR WE PROCEED TO S1
-- S8:  INTERRUPT STATE
-- FINISH:  STATE FOR COMING BACK TO FLOOR WITH LiftDir = 3


	-- instantiating the memory
	Memory0: entity work.MEMORY(RTL)
		port map (Address => Addr, Data => memory_data);

	-- instantiating the random_generator  
	RANDOM0: entity work.RANDOM_GENERATOR(RTL)
		port map (clk => clk, reset => reset, interrupt => interrupt, random_floor => random_floor);	
		

	 --%%%%%%%%%%%%%%%%%%%%% SEQUENTIAL SECTION %%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
	process (reset, clk)
	begin		
		if (reset = '1') then 
			pr_state <= S0; --go to S0
				
		elsif (clk'Event and clk = '1') then --in rising edge of the clock
			pr_state <= nx_state;  --go to next state
								
		end if;
		
	end process;
	
	
	--%%%%%%%%%%%%%%%%%%%%% NEXT STATE LOGIC %%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%	   
	process (pr_state, memory_data, start, count, interrupt)
	begin	
		
		
		--using case-when statements to determine the next state 
		case pr_state is 
				
			when S0 => 
				if (start = '1') then
					nx_state <= S1;					
				else 
					nx_state <= S0;					
				end if;
				
				
			when S1 =>
				nx_state <= S2;
		
				
			when S2 =>
				if (to_integer(unsigned(memory_data)) = 255) then
					-- Halt instruction (11111111)
					nx_state <= FINISH;
					
				else 
					nx_state <= S3;
					
				end if;
			
			when S3 =>
				nx_state <= S4;
				
				
			when S4 => 
				if (count = 0) then
					nx_state <= S5;	 
				else
					nx_state <= S4;
				end if;

			
			when S5 =>
				nx_state <= S6;
			
				
			when S6 => 
				if (count = 0) then
					nx_state <= S7;
				else
					nx_state <= S6;
				end if;
				
				
			
			when S7 =>
				if (interrupt = '1') then
					nx_state <= S8;
				else
					nx_state <= S1;
				end if;
					

				
			
			when S8 =>
				nx_state <= S3;
				
				
			when FINISH => 
				if (start = '1') then
					nx_state <= S1;
					
				else
					nx_state <= FINISH;
					
				end if;
				
				
				
			when others =>
				nx_state <= S0;
			
		end case;
		
	end process;
 
	
--%%%%%%%%%%%%%%%%%%%%% OUTPUT LOGIC %%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%

process (pr_state, memory_data)

-- The save variable is for saving the result of the multiplication and 
-- only assigning the 4 less significant bits.
variable save : std_logic_vector (7 downto 0);

-- for incrementing the address
variable inc : integer := 0;
begin 

	
	case pr_state is 
		
		when S0 =>
			Floor <= (others => '0');
			Timer <= (others => '0');
			LiftDir <= "00";
			LiftDoor <= '0';
			present_floor <= (others => '0'); -- ground floor 
			target_floor	  	 <= (others => '0'); 
			transition_time		 <= (others => '0');
			waiting_time 		 <= (others => '0');
			Addr <= (others => '0');
			inc := 0; 	
			
		when S1 =>
			target_floor <= memory_data (7 downto 4); -- fetching data from memory
			waiting_time <= memory_data (3 downto 0);
			Addr <= std_logic_vector(to_unsigned(inc, Addr'length));
		
		
		when S2 =>		
			
			-- transition time is the distance between two floors times 2 (2 secends for two adjacent floors)
			if (unsigned(target_floor) >= unsigned(present_floor)) then 
				save := std_logic_vector( ( unsigned(target_floor) - unsigned(present_floor) )  * 2 );
				transition_time <= save (3 downto 0);
			else 
				save := std_logic_vector( ( unsigned(present_floor) - unsigned(target_floor) )  * 2 );
				transition_time <= save (3 downto 0);
			end if;	

				
		
		when S3 =>	 
			inc := inc + 1;	 -- going to the next memory cell
			time_init <= to_integer(unsigned(transition_time));	-- time_init is transition_time
			
			
			
		
		when S4 =>
			Floor <= (others => '1'); -- transition state
			Timer <= (others => '0');
			LiftDoor <= '0';	
			if (target_floor > present_floor) then
				LiftDir <= "01"; -- going up
			else
				LiftDir <= "10"; -- going down
			end if;
			
			
			
		when S5 =>
			time_init <= to_integer(unsigned(waiting_time)); -- time_init is waiting_time
		   
			
		
		when S6 =>
			Floor <= target_floor; -- waiting state
			Timer <= std_logic_vector(to_unsigned(count, Timer'length));
			LiftDir <= "00";
			LiftDoor <= '1'; 
			present_floor <= target_floor;
			
		when S7 =>
			null; -- doing nothing
				
			
		when S8 =>	
			waiting_time <= "0101";	 -- 5 seconds
			target_floor <= random_floor;  -- the value from LFSR goes to target_floor
			LiftDoor <= '0';	 -- the door is closed
			
			
		when FINISH =>
			Floor <= (others => '0'); -- elevator is finished
			Timer <= (others => '0');
			LiftDir <= "11"; --waiting for the next list to come out
			LiftDoor <= '1';   -- the door is open
		
		
		when others => 
			Floor <= (others => '0');
			Timer <= (others => '0');
			LiftDir <= "00";
			LiftDoor <= '0';
			present_floor <= (others => '0');
		
			
	end case;
		
	
end process;



--%%%%%%%%%%%%%%%%%%%%% COUNTING PROCESS %%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
process (ONE_SECOND_CLOCK, pr_state, time_init)
variable time_count : integer := 0; 	 
variable s : integer := 0;
begin 
	
	-- This condition must run only one time when in S4 or S6
	if (s = 0) then
		time_count := time_init; 
		count <= time_count;
		s := 1;
	end if;
	
	-- This process is supposed to the the counting
	if ( pr_state = S4 or pr_state = S6 ) then
		
		if ( rising_edge(ONE_SECOND_CLOCK) ) then 
			time_count := time_count - 1; 
			count <= time_count;
		end if;
		

		
		
	else   
		-- This means the state is not S4 or S6 So we make s zero to initialize time_count with time_init
		s := 0;

	end if;	
	
	
	
end process;



	--%%%%%%%%%%%%%%%%%%%%% STATE DECODER %%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
	process (pr_state)
	begin  
		case pr_state is
			when S0 =>
				fsm_state <= "0000";	
			when S1 =>
				fsm_state <= "0001";
			when S2 =>
				fsm_state <= "0010";
			when S3 =>
				fsm_state <= "0011";
			when S4 =>
				fsm_state <= "0100";
			when S5 =>
				fsm_state <= "0101";
			when S6 =>
				fsm_state <= "0110";
			when S7 =>
				fsm_state <= "0111";	 
			when S8 =>
				fsm_state <= "1000";
			when finish =>
				fsm_state <= "1111";
			
			
			when others =>
			 	fsm_state <= "1010";
			
		end case;
		
	end process;  
	
	-- Showing middle signals in the simulation
	state <= fsm_state;	--putting the fsm_state signal into the port state 
	Memory_Out <= memory_data; --putting the memory_data signal inti the port Memory_Out  
	
	pres_floor <= present_floor;
	targ_floor <= target_floor;
	trans_time <= transition_time;
	wait_time <= waiting_time;
	address <= Addr;
	rand_floor <= random_floor;
	inter <= interrupt;
	counter_down <= count;
	time_initial <= time_init;


end architecture RTL;
